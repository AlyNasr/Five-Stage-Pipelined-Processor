LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
 
 
Entity Controlunit is 
port(
reset       :in std_logic;
opcode      :in std_logic_vector(4 downto 0);
C_Interrupt: in std_logic;

ALUop		:out std_logic_vector(3 downto 0);
ALUsrc		:out std_logic;
SpValue	:out std_logic_vector(2 downto 0);
   --Save		:out std_logic;
	 Restore	:out std_logic;
	 R1Data		:out std_logic_vector(1 downto 0);
	 RegDst		:out std_logic;
	 MemData	:out std_logic_vector(1 downto 0);
	 MemAddress	:out std_logic_vector(1 downto 0);
	 MemToReg	:out std_logic_vector(2 downto 0);
	 RegWrite1	:out std_logic;
	 RegWrite2	:out std_logic;
	 MemWrite	:out std_logic;
	 SetC		:out std_logic;
	 ClrC		:out std_logic;
	 JZ			:out std_logic;
	 JN			:out std_logic;
	 JC			:out std_logic;
	 JMP		:out std_logic;
	 Outp: out std_logic;
	 en_CCR: out std_logic;
	 Sp_en: out std_logic;
	 MemPc: out std_logic;
	 CF_en: out std_logic
	
);
end Controlunit;

ARCHITECTURE myControlUnit of Controlunit is
  Signal SMemWrite: std_logic;
  Signal Sen_CCR: std_logic;
  Signal SMemData: std_logic_vector(1 downto 0);
begin

process(reset,opcode)
  begin
    if (reset = '1') then
       ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			 Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			 SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ		<=	'0';
			 JN		<=	'0';
			 JC		<=	'0';
			 JMP		<=	'0';
			 Outp <= '0';
			 Sen_CCR <= '0';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '0';
   
   else
case opcode IS
when "00001" =>     -- setc
         ALUop		<=	"1100";
			   ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			R1Data		<=	"00";
			RegDst		<=	'0';
			SMemData		<=	"00";
			MemAddress	<=	"00";
			MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			SetC		<=	'1';
			ClrC		<=	'0';
			 JZ		<=	'0';
			 JN		<=	'0';
			 JC		<=	'0';
			 JMP		<=	'0';
			 Outp <= '0';
			 Sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
		-- ----	ClrC	----
		 when "00010" =>
			 ALUop		<=	"1011";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			MemAddress	<=	"00";
		  MemToReg	<= "000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'1';
			 JZ		<=	'0';
			 JN		<=	'0';
			 JC		<=	'0';
			 JMP		<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
-- ----	NOT		----
		 when "00011" =>
			 ALUop		<=	"1010";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
		  Restore		<=	'0';
			R1Data		<=	"10";
			 RegDst		<=	'0';
			 SMemData		<=	"00";
			MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '0'; 
-- ----	INC		----
		 when "00100" =>
			 ALUop		<=	"0001";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			 Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
		   ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
		-- ----	DEC		----
		 when "00101" =>
			 ALUop		<=	"0010";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<= "000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
			 -- ---		IN		----
		 when "00111" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			 SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"010";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ		<=	'0';
			 JN		<=	'0';
			 JC		<=	'0';
			 JMP		<=	'0';
			 Outp <= '0';
			 sen_CCR <= '0';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '0';
		-- ----	OUT		---
		 when "00110" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '1';
			 sen_CCR <= '0';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '0';
			-- ----	ADD		----
		 when "01001" =>
			 ALUop		<=	"0011";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
		-- ----	SUB		----
		when "01011" =>
			 ALUop		<=	"0101";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
		   Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
		-- ----	AND		----
		 when "01100" =>
			 ALUop		<=	"0110";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '0';
		-- ----	OR		----
		 when "01101" =>
			 ALUop		<=	"0111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
		   RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '0';
		-- ----	SWAP	----
		 when "01000" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"01";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"011";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'1';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '0';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '0';
		-- ----	AddI	----
		 when "01010" =>
			 ALUop		<=	"0011";
			 ALUsrc		<=	'1';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
		   Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
			 	-- ----	SHL		----
	 when "01110" =>
			 ALUop		<=	"1000";
			 ALUsrc		<=	'1';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
		-- ----	SHR		----
		 when "01111" =>
			 ALUop		<=	"1001";
			 ALUsrc		<=	'1';
			 SpValue		<=	"000";
			 --Save		<=	'0';
			 Restore		<=	'0';
			 R1Data		<=	"10";
			 RegDst		<=	'0';
			 SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
	     Outp <= '0';
			 sen_CCR <= '1';
			 Sp_en <= '0';
			 MemPc <= '0';
			 CF_en <= '1';
			 -- ----	PUSH	----
		 when "10000" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"001";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"01";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'1';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '0';
			 Sp_en <= '1';
	     MemPc <= '0';
	     CF_en <= '0';
		-- ----	POP		----
		 when "10001" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"010";
			-- Save		<=	'0';
			 Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"01";
			 MemToReg	<=	"001";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '0';
			 Sp_en <= '1';
	     MemPc <= '0';
	     CF_en <= '0';
		-- ----	LDM		----
		 when "10010" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"111";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '0';
			 Sp_en <= '0';
	     MemPc <= '0';
	     CF_en <= '0';
		-- ----	LDD		----
		 when "10011" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			 Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"10";
			 MemToReg	<=	"001";
			 RegWrite1	<=	'1';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			sen_CCR <= '0';
	     Sp_en <= '0';
	     MemPc <= '0';
	     CF_en <= '0';
		-- ----	STD		----
		 when "10100" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"10";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'1';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
       Outp <= '0';
			 sen_CCR <= '0';
	     Sp_en <= '0';
	     MemPc <= '0';
	     CF_en <= '0';
	 -- ----	JZ		----
		 when "10101" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'1';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
	     Sp_en <= '0';
	     MemPc <= '0';
	     CF_en <= '0';
		-- ----	JN		----
		 when "10110" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'1';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
	     Sp_en <= '0';
       MemPc <= '0';
       CF_en <= '0';
		-- ----	JC		----	
		 when "10111" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'1';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
	     Sp_en <= '0';
       MemPc <= '0';
       CF_en <= '0';
		-- ----	JMP		----
		 when "11000" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
			 Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			JMP			<=	'1';
			   Outp <= '0';
			   sen_CCR <= '0';
	       Sp_en <= '0';
         MemPc <= '0';
         CF_en <= '0';
		-- ----	RET		----
	 when "11010" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"100";
			-- Save		<=	'0';
			 Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			 SMemData		<=	"00";
			 MemAddress	<=	"01";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 SMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '0';
	     Sp_en <= '1';
       MemPc <= '1';
       CF_en <= '0';
		-- ----	RTI		----
		 when "11011" =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"011";
			-- Save		<=	'0';
			 Restore		<=	'1';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			 SMemData		<=	"00";
			 MemAddress	<=	"01";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 SMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '1';
	     Sp_en <= '1';
       MemPc <= '1';
       CF_en <= '0';
		-- ----	CALL	----
		 when "11001" =>
		 ALUop		<=	"1111";
		 ALUsrc		<=	'0';
			 SpValue		<=	"110";
			-- Save		<=	'0';
			 Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			 SMemData		<=	"10";
			 MemAddress	<=	"01";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 SMemWrite	<=	'1';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'1';
		   Outp <= '0';
			 sen_CCR <= '0';
	     Sp_en <= '1';
       MemPc <= '0';
       CF_en <= '0';
		 when others =>
			 ALUop		<=	"1111";
			 ALUsrc		<=	'0';
			 SpValue		<=	"000";
			-- Save		<=	'0';
		   Restore		<=	'0';
			 R1Data		<=	"00";
			 RegDst		<=	'0';
			 SMemData		<=	"00";
			 MemAddress	<=	"00";
			 MemToReg	<=	"000";
			 RegWrite1	<=	'0';
			 RegWrite2	<=	'0';
			 sMemWrite	<=	'0';
			 SetC		<=	'0';
			 ClrC		<=	'0';
			 JZ			<=	'0';
			 JN			<=	'0';
			 JC			<=	'0';
			 JMP			<=	'0';
			 Outp <= '0';
			 sen_CCR <= '0';
       Sp_en <= '0';
       MemPc <= '0';
       CF_en <= '0';
   end case;
  end if;
end process;
 MemWrite <= '1' WHEN C_Interrupt = '1'
        ELSE sMemWrite;
 en_CCR <= '1' WHEN C_Interrupt = '1'
      ELSE   sen_CCR ; 
 MemData <= "01" WHEN C_Interrupt = '1'
      Else SMemData;            
End myControlUnit;
